module SPI_mnrch (
    input logic clk,            // System clock driving the controller
    input logic rst_n,          // Active-low asynchronous reset
    input logic MISO,           // Master-In-Slave-Out (data from slave)
    input logic wrt,            // Start transfer request (one-shot or level)
    input logic [15:0] wt_data, // 16-bit data to transmit (MSB first)
    output logic MOSI,          // Master-Out-Slave-In (data to slave)
    output logic SCLK,          // SPI serial clock (generated by this module)
    output logic SS_n,          // Active-low slave select (chip select)
    output logic done,          // Pulse/level signaling transfer completion
    output logic [15:0] rd_data // 16-bit data received from slave
);

logic [3:0] SCLK_div;           // 4-bit clock divider/counter for SCLK generation (clk/16)
logic ld_SCLK, smpl, MISO_smpl, init, set_done, done15, shft_im, shft;
logic [15:0] shft_reg;          // Shift register for TX (MOSI) and RX (MISO) data
logic [3:0] bit_cnt;            // Counts number of bits shifted (0..15)



always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        SCLK_div <= 4'b1011;   // Reset SCLK divider to a known phase
    end else if (ld_SCLK) begin
        SCLK_div <= 4'b1011;   // Reload to align SCLK phase for next transaction
    end else begin
        SCLK_div <= SCLK_div + 4'd1; // Free-run increment
    end
end

assign SCLK = SCLK_div[3];          // SCLK toggles every 8 cycles of 'clk' (50% duty)
assign smpl = (SCLK_div == 4'b0111); // Sample point relative to SCLK low-high boundary
assign shft_im = (SCLK_div == 4'b1111); // Shift point near the high-low boundary


always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n)          
     MISO_smpl <= 1'b0;        // Default captured value on reset
  else if (smpl)        
    MISO_smpl <= MISO;         // Sample MISO at defined divider tap
end

always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        shft_reg <= 16'd0;     // Clear on reset
    end
    else if (init) begin
        shft_reg <= wt_data;    // Load data to transmit
    end
    else if (shft) begin
        shft_reg <= {shft_reg[14:0], MISO_smpl}; // Shift out MSB, shift in sampled MISO
    end
end
assign MOSI = shft_reg[15];     // Drive MOSI with current MSB (MSB-first protocol)
assign rd_data = shft_reg;      // Expose received/shifted data to output


always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        bit_cnt <= 4'd0;
    end
    else if (init) begin
        bit_cnt <= 4'd0;        // Prepare to count a new 16-bit transfer
    end
    else if (shft) begin
        bit_cnt <= bit_cnt + 4'd1; // Count each shift event
    end
    else begin
        bit_cnt <= bit_cnt;     // Hold
    end
end

assign done15 = &bit_cnt;       // High when bit_cnt == 4'b1111 (15)

// FSM encoding for transaction control
typedef enum logic [1:0] {
    IDLE,       
    TRANSFER,    
    COMPLETE,    
    FRONTPORCH   
} state_t;

state_t state, nxt_state;

// State register
always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        state <= IDLE;
    end else begin
        state <= nxt_state;
    end
end

always_comb begin
    // Default assignments
    ld_SCLK = 1'b1;    // Hold divider unless actively transferring
    init = 1'b0;
    set_done = 1'b0;
    nxt_state = state;
    shft = 1'b0;

    case (state)
        IDLE: begin
            if (wrt) begin
                ld_SCLK = 1'b0; // Release divider to start SCLK
                init = 1'b1;    // Load shift register and assert SS_n
                nxt_state = FRONTPORCH; // Allow phase to settle before first shift
            end
        end
    FRONTPORCH: begin
        ld_SCLK = 1'b0;         // Keep SCLK running
        if (shft_im) begin
            nxt_state = TRANSFER; // Enter shifting on specific divider tap
        end else begin
            nxt_state = FRONTPORCH;
        end
    end
        TRANSFER: begin 
        ld_SCLK = 1'b0;         // Keep SCLK running during transfer
        if (done15) begin        // After 15 shifts, move to COMPLETE for final shift
            nxt_state = COMPLETE;
        end else begin
            if (shft_im) begin
                shft = 1'b1;    // Shift once per SCLK period at the defined tap
            end
            nxt_state = TRANSFER;
            end
        end
        COMPLETE: begin
            ld_SCLK = 1'b0;     // Keep SCLK active until final shift occurs
            if (shft_im) begin
                shft = 1'b1;    // Perform the 16th and final shift
                set_done = 1'b1; // Flag completion and end the transaction
                ld_SCLK = 1'b1; // Reload divider to stop/realign SCLK post-transfer
                nxt_state = IDLE;
            end else
                nxt_state = COMPLETE;
        end
    endcase
end

always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        SS_n <= 1'b1;           // Inactive (no slave selected) on reset
    end else if (init) begin
        SS_n <= 1'b0;           // Select slave at start of transfer
    end
    else if (set_done) begin
        SS_n <= 1'b1;           // Release slave at end of transfer
    end
end

always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        done <= 1'b0;
    end else if (set_done) begin
        done <= 1'b1;
    end else if (init) begin
        done <= 1'b0;
    end
end



endmodule